<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-18.6623,-46.7485,68.4042,-124.348</PageViewport>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW</type>
<position>1,-69.5</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>4 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>1,-82.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>5 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_DFF_LOW</type>
<position>1,-95.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-12,-64.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_NAND2</type>
<position>14,-76.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>9,-77.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>BA_NAND2</type>
<position>14,-89.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>9,-90.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>19,-76.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>19,-89.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AE_DFF_LOW</type>
<position>1,-108.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>14,-102.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AE_SMALL_INVERTER</type>
<position>9,-103.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>19,-102.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND2</type>
<position>14,-115.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_SMALL_INVERTER</type>
<position>9,-116.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>19,-115.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>-12,-59.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>-3,-60.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_DFF_LOW</type>
<position>37,-71</position>
<input>
<ID>IN_0</ID>105 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_DFF_LOW</type>
<position>37,-84</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>37,-97</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>24,-66</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>BA_NAND2</type>
<position>50,-78</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>45,-79</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>BA_NAND2</type>
<position>50,-91</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_SMALL_INVERTER</type>
<position>45,-92</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>55,-78</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>55,-91</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>37,-110</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>80 </output>
<input>
<ID>clock</ID>66 </input>
<gparam>angle 270</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_NAND2</type>
<position>50,-104</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_SMALL_INVERTER</type>
<position>45,-105</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>55,-104</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>BA_NAND2</type>
<position>50,-117</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>45,-118</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>55,-117</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>24,-61</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_OR2</type>
<position>33,-62</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_AND2</type>
<position>39,-65</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_TOGGLE</type>
<position>24,-56</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-116.5,-5,-64.5</points>
<intersection>-116.5 26</intersection>
<intersection>-103.5 20</intersection>
<intersection>-90.5 6</intersection>
<intersection>-77.5 3</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-64.5,1.09512e-007,-64.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-5 0</intersection>
<intersection>1.09512e-007 30</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-5,-77.5,7,-77.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection>
<intersection>1.09512e-007 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-5,-90.5,7,-90.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection>
<intersection>1.09512e-007 22</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1.09512e-007,-79.5,1.09512e-007,-77.5</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>-77.5 3</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-5,-103.5,7,-103.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection>
<intersection>1.09512e-007 29</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>1.09512e-007,-92.5,1.09512e-007,-90.5</points>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<intersection>-90.5 6</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-5,-116.5,7,-116.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>1.09512e-007,-105.5,1.09512e-007,-103.5</points>
<connection>
<GID>11</GID>
<name>clock</name></connection>
<intersection>-103.5 20</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>1.09512e-007,-66.5,1.09512e-007,-64.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>-64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-77.5,11,-77.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-90.5,11,-90.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-79.5,3,-72.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>3,-75.5,11,-75.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-92.5,3,-85.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-88.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>3,-88.5,11,-88.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>17,-76.5,18,-76.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>9</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>17,-89.5,18,-89.5</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-103.5,11,-103.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-105.5,3,-98.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-101.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>3,-101.5,11,-101.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>17,-102.5,18,-102.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-116.5,11,-116.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-114.5,-7,-61.5</points>
<intersection>-114.5 3</intersection>
<intersection>-61.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-7,-114.5,11,-114.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection>
<intersection>3 8</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-7,-61.5,-6,-61.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-7 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>3,-114.5,3,-111.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-114.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>17,-115.5,18,-115.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-59.5,-6,-59.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-66.5,3,-60.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-60.5,3,-60.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-118,31,-66</points>
<intersection>-118 26</intersection>
<intersection>-105 20</intersection>
<intersection>-92 6</intersection>
<intersection>-79 3</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-66,36,-66</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection>
<intersection>36 30</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-79,43,-79</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection>
<intersection>36 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>31,-92,43,-92</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection>
<intersection>36 22</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>36,-81,36,-79</points>
<connection>
<GID>77</GID>
<name>clock</name></connection>
<intersection>-79 3</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>31,-105,43,-105</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection>
<intersection>36 29</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>36,-94,36,-92</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>-92 6</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>31,-118,43,-118</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>36,-107,36,-105</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>-105 20</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>36,-68,36,-66</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-79,47,-79</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-92,47,-92</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-81,39,-74</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-77 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>39,-77,47,-77</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-94,39,-87</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-90 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>39,-90,47,-90</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>53,-78,54,-78</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<connection>
<GID>82</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>53,-91,54,-91</points>
<connection>
<GID>92</GID>
<name>N_in0</name></connection>
<connection>
<GID>85</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-105,47,-105</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-107,39,-100</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-103 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>39,-103,47,-103</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>53,-104,54,-104</points>
<connection>
<GID>100</GID>
<name>N_in0</name></connection>
<connection>
<GID>98</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-118,47,-118</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-116,29,-63</points>
<intersection>-116 3</intersection>
<intersection>-63 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>29,-116,47,-116</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection>
<intersection>39 8</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>29,-63,30,-63</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>39,-116,39,-113</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-116 3</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>53,-117,54,-117</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>104</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-61,30,-61</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-68,39,-68</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-62,38,-62</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-62,40,-56</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-56,40,-56</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 1>
<page 2>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 2>
<page 3>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 3>
<page 4>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 4>
<page 5>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 5>
<page 6>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 6>
<page 7>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 7>
<page 8>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 8>
<page 9>
<PageViewport>-17.75,0,47.55,-58.2</PageViewport></page 9></circuit>